library ieee;
use ieee.std_logic_1164.all;

entity memory_state_machine is

	port(
		clk		 	: in	std_logic;
		ReqLeit	 	: inout	std_logic;
		Ack			: inout	std_logic;
		reset	 	: in	std_logic;
		output	 	: out	std_logic_vector(1 downto 0)
	);

end entity;

architecture rtl of memory_state_machine is

	-- Build an enumerated type for the state machine
	type state_type is (s0, s1, s2, s3);

	-- Register to hold the current state
	signal state : state_type;

begin

	process (clk, reset) begin

		if reset = '1' then
			state <= s0;

		elsif (rising_edge(clk)) then

			-- Determine the next state synchronously, based on
			-- the current state and the input
			case state is
				when s0=>
					if ReqLeit = '1' then
						state <= s1;
					else
						state <= s0;
					end if;
				when s1=>
					if ReqLeit = '1' then
						state <= s2;
					else
						state <= s1;
					end if;
				when s2=>
					if ReqLeit = '1' then
						state <= s3;
					else
						state <= s2;
					end if;
				when s3=>
					if ReqLeit = '1' then
						state <= s3;
					else
						state <= s1;
					end if;
			end case;

		end if;
	end process;

	-- Determine the output based only on the current state
	-- and the input (do not wait for a clock edge).
	process (state, ReqLeit)
	begin
			case state is
				when s0=>
					if ReqLeit = '1' then
						output <= "00";
					else
						output <= "01";
					end if;
				when s1=>
					if ReqLeit = '1' then
						output <= "01";
					else
						output <= "11";
					end if;
				when s2=>
					if ReqLeit = '1' then
						output <= "10";
					else
						output <= "10";
					end if;
				when s3=>
					if ReqLeit = '1' then
						output <= "11";
					else
						output <= "10";
					end if;
			end case;
	end process;

end rtl;
